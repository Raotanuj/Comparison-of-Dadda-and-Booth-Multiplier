module Dadda (A, B, Mul);

parameter N = 16;

input [N-1:0] A, B;
output [2*N-1:0] Mul;

wire S2[31:0][15:0];
//reg S3[8:0][8:0];
//wire S3[31:9][15:0];
wire S3[31:0][15:0];
wire S4[31:0][15:0];
wire S5[31:0][15:0];
wire S6[31:0][15:0];
wire S7[31:0][15:0];

reg S1[15:0][15:0];

integer i,j;

always @(*) begin			// Initialize the partial products

	for(i=0;i<N;i=i+1) begin

		for(j=0;j<N;j=j+1) begin
	
			S1[i][j] = A[i] & B[j];
		end
	end
end


// S1 - Stage-1 

assign S2[0][0] = S1[0][0];

assign S2[1][0] = S1[1][0];
assign S2[1][1] = S1[0][1];

assign S2[2][0] = S1[2][0];
assign S2[2][1] = S1[1][1];
assign S2[2][2] = S1[0][2];

assign S2[3][0] = S1[3][0];
assign S2[3][1] = S1[2][1];
assign S2[3][2] = S1[1][2];
assign S2[3][3] = S1[0][3];

assign S2[4][0] = S1[4][0];
assign S2[4][1] = S1[3][1];
assign S2[4][2] = S1[2][2];
assign S2[4][3] = S1[1][3];
assign S2[4][4] = S1[0][4];

assign S2[5][0] = S1[5][0];
assign S2[5][1] = S1[4][1];
assign S2[5][2] = S1[3][2];
assign S2[5][3] = S1[2][3];
assign S2[5][4] = S1[1][4];
assign S2[5][5] = S1[0][5];

assign S2[6][0] = S1[6][0];
assign S2[6][1] = S1[5][1];
assign S2[6][2] = S1[4][2];
assign S2[6][3] = S1[3][3];
assign S2[6][4] = S1[2][4];
assign S2[6][5] = S1[1][5];
assign S2[6][6] = S1[0][6];

assign S2[7][0] = S1[7][0];
assign S2[7][1] = S1[6][1];
assign S2[7][2] = S1[5][2];
assign S2[7][3] = S1[4][3];
assign S2[7][4] = S1[3][4];
assign S2[7][5] = S1[2][5];
assign S2[7][6] = S1[1][6];
assign S2[7][7] = S1[0][7];

assign S2[8][0] = S1[8][0];
assign S2[8][1] = S1[7][1];
assign S2[8][2] = S1[6][2];
assign S2[8][3] = S1[5][3];
assign S2[8][4] = S1[4][4];
assign S2[8][5] = S1[3][5];
assign S2[8][6] = S1[2][6];
assign S2[8][7] = S1[1][7];
assign S2[8][8] = S1[0][8];

assign S2[9][0] = S1[9][0];
assign S2[9][1] = S1[8][1];
assign S2[9][2] = S1[7][2];
assign S2[9][3] = S1[6][3];
assign S2[9][4] = S1[5][4];
assign S2[9][5] = S1[4][5];
assign S2[9][6] = S1[3][6];
assign S2[9][7] = S1[2][7];
assign S2[9][8] = S1[1][8];
assign S2[9][9] = S1[0][9];

assign S2[10][0] = S1[10][0];
assign S2[10][1] = S1[9][1];
assign S2[10][2] = S1[8][2];
assign S2[10][3] = S1[7][3];
assign S2[10][4] = S1[6][4];
assign S2[10][5] = S1[5][5];
assign S2[10][6] = S1[4][6];
assign S2[10][7] = S1[3][7];
assign S2[10][8] = S1[2][8];
assign S2[10][9] = S1[1][9];
assign S2[10][10] = S1[0][10];

assign S2[11][0] = S1[11][0];
assign S2[11][1] = S1[10][1];
assign S2[11][2] = S1[9][2];
assign S2[11][3] = S1[8][3];
assign S2[11][4] = S1[7][4];
assign S2[11][5] = S1[6][5];
assign S2[11][6] = S1[5][6];
assign S2[11][7] = S1[4][7];
assign S2[11][8] = S1[3][8];
assign S2[11][9] = S1[2][9];
assign S2[11][10] = S1[1][10];
assign S2[11][11] = S1[0][11];

HA H1 (S1[12][0], S1[11][1], S2[12][0], S2[13][0]);
assign S2[12][1] = S1[10][2];
assign S2[12][2] = S1[9][3];
assign S2[12][3] = S1[8][4];
assign S2[12][4] = S1[7][5];
assign S2[12][5] = S1[6][6];
assign S2[12][6] = S1[5][7];
assign S2[12][7] = S1[4][8];
assign S2[12][8] = S1[3][9];
assign S2[12][9] = S1[2][10];
assign S2[12][10] = S1[1][11];
assign S2[12][11] = S1[0][12];

FA F1 (S1[13][0], S1[12][1], S1[11][2], S2[13][1], S2[14][0]);
HA H2 (S1[10][3], S1[9][4], S2[13][2], S2[14][1]);
assign S2[13][3] = S1[8][5];
assign S2[13][4] = S1[7][6];
assign S2[13][5] = S1[6][7];
assign S2[13][6] = S1[5][8];
assign S2[13][7] = S1[4][9];
assign S2[13][8] = S1[3][10];
assign S2[13][9] = S1[2][11];
assign S2[13][10] = S1[1][12];
assign S2[13][11] = S1[0][13];

FA F2 (S1[14][0], S1[13][1], S1[12][2], S2[14][2], S2[15][0]);
FA F3 (S1[11][3], S1[10][4], S1[9][5], S2[14][3], S2[15][1]);
HA H3 (S1[8][6], S1[7][7], S2[14][4], S2[15][2]);
assign S2[14][5] = S1[6][8];
assign S2[14][6] = S1[5][9];
assign S2[14][7] = S1[4][10];
assign S2[14][8] = S1[3][11];
assign S2[14][9] = S1[2][12];
assign S2[14][10] = S1[1][13];
assign S2[14][11] = S1[0][14];

FA F4 (S1[15][0], S1[14][1], S1[13][2], S2[15][3], S2[16][0]);
FA F5 (S1[12][3], S1[11][4], S1[10][5], S2[15][4], S2[16][1]);
FA F6 (S1[9][6], S1[8][7], S1[7][8], S2[15][5], S2[16][2]);
HA H4 (S1[6][9], S1[5][10], S2[15][6], S2[16][3]);
assign S2[15][7] = S1[4][11];
assign S2[15][8] = S1[3][12];
assign S2[15][9] = S1[2][13];
assign S2[15][10] = S1[1][14];
assign S2[15][11] = S1[0][15];

FA F14 (S1[15][1], S1[14][2], S1[13][3], S2[16][4], S2[17][0]);
FA F15 (S1[12][4], S1[11][5], S1[10][6], S2[16][5], S2[17][1]);
FA F7 (S1[9][7], S1[8][8], S1[7][9], S2[16][6], S2[17][2]);
HA H5 (S1[6][10], S1[5][11], S2[16][7], S2[17][3]);
assign S2[16][8] = S1[4][12];
assign S2[16][9] = S1[3][13];
assign S2[16][10] = S1[2][14];
assign S2[16][11] = S1[1][15];

FA F8  (S1[15][2], S1[14][3], S1[13][4], S2[17][4], S2[18][0]);
FA F9  (S1[12][5], S1[11][6], S1[10][7], S2[17][5], S2[18][1]);
FA F10 (S1[9][8], S1[8][9], S1[7][10], S2[17][6], S2[18][2]);
assign S2[17][7] = S1[6][11];
assign S2[17][8] = S1[5][12];
assign S2[17][9] = S1[4][13];
assign S2[17][10] = S1[3][14];
assign S2[17][11] = S1[2][15];

FA F11 (S1[15][3], S1[14][4], S1[13][5], S2[18][3], S2[19][0]);
FA F12 (S1[12][6], S1[11][7], S1[10][8], S2[18][4], S2[19][1]);
assign S2[18][5] = S1[9][9];
assign S2[18][6] = S1[8][10];
assign S2[18][7] = S1[7][11];
assign S2[18][8] = S1[6][12];
assign S2[18][9] = S1[5][13];
assign S2[18][10] = S1[4][14];
assign S2[18][11] = S1[3][15];

FA F13 (S1[15][4], S1[14][5], S1[13][6], S2[19][2], S2[20][0]);
assign S2[19][3] = S1[12][7];
assign S2[19][4] = S1[11][8];
assign S2[19][5] = S1[10][9];
assign S2[19][6] = S1[9][10];
assign S2[19][7] = S1[8][11];
assign S2[19][8] = S1[7][12];
assign S2[19][9] = S1[6][13];
assign S2[19][10] = S1[5][14];
assign S2[19][11] = S1[4][15];

assign S2[20][1] = S1[15][5];
assign S2[20][2] = S1[14][6];
assign S2[20][3] = S1[13][7];
assign S2[20][4] = S1[12][8];
assign S2[20][5] = S1[11][9];
assign S2[20][6] = S1[10][10];
assign S2[20][7] = S1[9][11];
assign S2[20][8] = S1[8][12];
assign S2[20][9] = S1[7][13];
assign S2[20][10] = S1[6][14];
assign S2[20][11] = S1[5][15];

assign S2[21][0] = S1[15][6];
assign S2[21][1] = S1[14][7];
assign S2[21][2] = S1[13][8];
assign S2[21][3] = S1[12][9];
assign S2[21][4] = S1[11][10];
assign S2[21][5] = S1[10][11];
assign S2[21][6] = S1[9][12];
assign S2[21][7] = S1[8][13];
assign S2[21][8] = S1[7][14];
assign S2[21][9] = S1[6][15];

assign S2[22][0] = S1[15][7];
assign S2[22][1] = S1[14][8];
assign S2[22][2] = S1[13][9];
assign S2[22][3] = S1[12][10];
assign S2[22][4] = S1[11][11];
assign S2[22][5] = S1[10][12];
assign S2[22][6] = S1[9][13];
assign S2[22][7] = S1[8][14];
assign S2[22][8] = S1[7][15];

assign S2[23][0] = S1[15][8];
assign S2[23][1] = S1[14][9];
assign S2[23][2] = S1[13][10];
assign S2[23][3] = S1[12][11];
assign S2[23][4] = S1[11][12];
assign S2[23][5] = S1[10][13];
assign S2[23][6] = S1[9][14];
assign S2[23][7] = S1[8][15];

assign S2[24][0] = S1[15][9];
assign S2[24][1] = S1[14][10];
assign S2[24][2] = S1[13][11];
assign S2[24][3] = S1[12][12];
assign S2[24][4] = S1[11][13];
assign S2[24][5] = S1[10][14];
assign S2[24][6] = S1[9][15];

assign S2[25][0] = S1[15][10];
assign S2[25][1] = S1[14][11];
assign S2[25][2] = S1[13][12];
assign S2[25][3] = S1[12][13];
assign S2[25][4] = S1[11][14];
assign S2[25][5] = S1[10][15];

assign S2[26][0] = S1[15][11];
assign S2[26][1] = S1[14][12];
assign S2[26][2] = S1[13][13];
assign S2[26][3] = S1[12][14];
assign S2[26][4] = S1[11][15];

assign S2[27][0] = S1[15][12];
assign S2[27][1] = S1[14][13];
assign S2[27][2] = S1[13][14];
assign S2[27][3] = S1[12][15];

assign S2[28][0] = S1[15][13];
assign S2[28][1] = S1[14][14];
assign S2[28][2] = S1[13][15];

assign S2[29][0] = S1[15][14];
assign S2[29][1] = S1[14][15];

assign S2[30][0] = S1[15][15];



// S2 - Stage-2 			


 assign S3[0][0] = S2[0][0];

 assign S3[1][0] = S2[1][0];
 assign S3[1][1] = S2[1][1];

 assign S3[2][0] = S2[2][0];
 assign S3[2][1] = S2[2][1];
 assign S3[2][2] = S2[2][2];

 assign S3[3][0] = S2[3][0];
 assign S3[3][1] = S2[3][1];
 assign S3[3][2] = S2[3][2];
 assign S3[3][3] = S2[3][3];

 assign S3[4][0] = S2[4][0];
 assign S3[4][1] = S2[4][1];
 assign S3[4][2] = S2[4][2];
 assign S3[4][3] = S2[4][3];
 assign S3[4][4] = S2[4][4];

 assign S3[5][0] = S2[5][0];
 assign S3[5][1] = S2[5][1];
 assign S3[5][2] = S2[5][2];
 assign S3[5][3] = S2[5][3];
 assign S3[5][4] = S2[5][4];
 assign S3[5][5] = S2[5][5];

 assign S3[6][0] = S2[6][0];
 assign S3[6][1] = S2[6][1];
 assign S3[6][2] = S2[6][2];
 assign S3[6][3] = S2[6][3];
 assign S3[6][4] = S2[6][4];
 assign S3[6][5] = S2[6][5];
 assign S3[6][6] = S2[6][6];

 assign S3[7][0] = S2[7][0];
 assign S3[7][1] = S2[7][1];
 assign S3[7][2] = S2[7][2];
 assign S3[7][3] = S2[7][3];
 assign S3[7][4] = S2[7][4];
 assign S3[7][5] = S2[7][5];
 assign S3[7][6] = S2[7][6];
 assign S3[7][7] = S2[7][7];

 assign S3[8][0] = S2[8][0];
 assign S3[8][1] = S2[8][1];
 assign S3[8][2] = S2[8][2];
 assign S3[8][3] = S2[8][3];
 assign S3[8][4] = S2[8][4];
 assign S3[8][5] = S2[8][5];
 assign S3[8][6] = S2[8][6];
 assign S3[8][7] = S2[8][7];
 assign S3[8][8] = S2[8][8];



HA H201 (S2[9][0], S2[9][1], S3[9][0], S3[10][0]);
assign S3[9][1] = S2[9][2];
assign S3[9][2] = S2[9][3];
assign S3[9][3] = S2[9][4];
assign S3[9][4] = S2[9][5];
assign S3[9][5] = S2[9][6];
assign S3[9][6] = S2[9][7];
assign S3[9][7] = S2[9][8];
assign S3[9][8] = S2[9][9];

FA F201 (S2[10][0], S2[10][1], S2[10][2], S3[10][1], S3[11][0]);
HA H202 (S2[10][3], S2[10][4], S3[10][2], S3[11][1]);
assign S3[10][3] = S2[10][5];
assign S3[10][4] = S2[10][6];
assign S3[10][5] = S2[10][7];
assign S3[10][6] = S2[10][8];
assign S3[10][7] = S2[10][9];
assign S3[10][8] = S2[10][10];

FA F202 (S2[11][0], S2[11][1], S2[11][2], S3[11][2], S3[12][0]);
FA F203 (S2[11][3], S2[11][4], S2[11][5], S3[11][3], S3[12][1]);
HA H203 (S2[11][6], S2[11][7], S3[11][4], S3[12][2]);
assign S3[11][5] = S2[11][8];
assign S3[11][6] = S2[11][9];
assign S3[11][7] = S2[11][10];
assign S3[11][8] = S2[11][11];

FA F204 (S2[12][0], S2[12][1], S2[12][2], S3[12][3], S3[13][0]);
FA F205 (S2[12][3], S2[12][4], S2[12][5], S3[12][4], S3[13][1]);
FA F206 (S2[12][6], S2[12][7], S2[12][8], S3[12][5], S3[13][2]);
assign S3[12][6] = S2[12][9];
assign S3[12][7] = S2[12][10];
assign S3[12][8] = S2[12][11];

FA F207 (S2[13][0], S2[13][1], S2[13][2], S3[13][3], S3[14][0]);
FA F208 (S2[13][3], S2[13][4], S2[13][5], S3[13][4], S3[14][1]);
FA F209 (S2[13][6], S2[13][7], S2[13][8], S3[13][5], S3[14][2]);
assign S3[13][6] = S2[13][9];
assign S3[13][7] = S2[13][10];
assign S3[13][8] = S2[13][11];

FA F210 (S2[14][0], S2[14][1], S2[14][2], S3[14][3], S3[15][0]);
FA F211 (S2[14][3], S2[14][4], S2[14][5], S3[14][4], S3[15][1]);
FA F212 (S2[14][6], S2[14][7], S2[14][8], S3[14][5], S3[15][2]);
assign S3[14][6] = S2[14][9];
assign S3[14][7] = S2[14][10];
assign S3[14][8] = S2[14][11];

FA F213 (S2[15][0], S2[15][1], S2[15][2], S3[15][3], S3[16][0]);
FA F214 (S2[15][3], S2[15][4], S2[15][5], S3[15][4], S3[16][1]);
FA F215 (S2[15][6], S2[15][7], S2[15][8], S3[15][5], S3[16][2]);
assign S3[15][6] = S2[15][9];
assign S3[15][7] = S2[15][10];
assign S3[15][8] = S2[15][11];

FA F216 (S2[16][0], S2[16][1], S2[16][2], S3[16][3], S3[17][0]);
FA F217 (S2[16][3], S2[16][4], S2[16][5], S3[16][4], S3[17][1]);
FA F218 (S2[16][6], S2[16][7], S2[16][8], S3[16][5], S3[17][2]);
assign S3[16][6] = S2[16][9];
assign S3[16][7] = S2[16][10];
assign S3[16][8] = S2[16][11];

FA F219 (S2[17][0], S2[17][1], S2[17][2], S3[17][3], S3[18][0]);
FA F220 (S2[17][3], S2[17][4], S2[17][5], S3[17][4], S3[18][1]);
FA F221 (S2[17][6], S2[17][7], S2[17][8], S3[17][5], S3[18][2]);
assign S3[17][6] = S2[17][9];
assign S3[17][7] = S2[17][10];
assign S3[17][8] = S2[17][11];

FA F222 (S2[18][0], S2[18][1], S2[18][2], S3[18][3], S3[19][0]);
FA F223 (S2[18][3], S2[18][4], S2[18][5], S3[18][4], S3[19][1]);
FA F224 (S2[18][6], S2[18][7], S2[18][8], S3[18][5], S3[19][2]);
assign S3[18][6] = S2[18][9];
assign S3[18][7] = S2[18][10];
assign S3[18][8] = S2[18][11];

FA F225 (S2[19][0], S2[19][1], S2[19][2], S3[19][3], S3[20][0]);
FA F226 (S2[19][3], S2[19][4], S2[19][5], S3[19][4], S3[20][1]);
FA F227 (S2[19][6], S2[19][7], S2[19][8], S3[19][5], S3[20][2]);
assign S3[19][6] = S2[19][9];
assign S3[19][7] = S2[19][10];
assign S3[19][8] = S2[19][11];

FA F228 (S2[20][0], S2[20][1], S2[20][2], S3[20][3], S3[21][0]);
FA F229 (S2[20][3], S2[20][4], S2[20][5], S3[20][4], S3[21][1]);
FA F230 (S2[20][6], S2[20][7], S2[20][8], S3[20][5], S3[21][2]);
assign S3[20][6] = S2[20][9];
assign S3[20][7] = S2[20][10];
assign S3[20][8] = S2[20][11];


FA F231 (S2[21][0], S2[21][1], S2[21][2], S3[21][3], S3[22][0]);
FA F232 (S2[21][3], S2[21][4], S2[21][5], S3[21][4], S3[22][1]);
assign S3[21][5] = S2[21][6];
assign S3[21][6] = S2[21][7];
assign S3[21][7] = S2[21][8];
assign S3[21][8] = S2[21][9];

FA F233 (S2[22][0], S2[22][1], S2[22][2], S3[22][2], S3[23][0]);
assign S3[22][3] = S2[22][3];
assign S3[22][4] = S2[22][4];
assign S3[22][5] = S2[22][5];
assign S3[22][6] = S2[22][6];
assign S3[22][7] = S2[22][7];
assign S3[22][8] = S2[22][8];

assign S3[23][1] = S2[23][0];
assign S3[23][2] = S2[23][1];
assign S3[23][3] = S2[23][2];
assign S3[23][4] = S2[23][3];
assign S3[23][5] = S2[23][4];
assign S3[23][6] = S2[23][5];
assign S3[23][7] = S2[23][6];
assign S3[23][8] = S2[23][7];

assign S3[24][0] = S2[24][0];
assign S3[24][1] = S2[24][1];
assign S3[24][2] = S2[24][2];
assign S3[24][3] = S2[24][3];
assign S3[24][4] = S2[24][4];
assign S3[24][5] = S2[24][5];
assign S3[24][6] = S2[24][6];

assign S3[25][0] = S2[25][0];
assign S3[25][1] = S2[25][1];
assign S3[25][2] = S2[25][2];
assign S3[25][3] = S2[25][3];
assign S3[25][4] = S2[25][4];
assign S3[25][5] = S2[25][5];

assign S3[26][0] = S2[26][0];
assign S3[26][1] = S2[26][1];
assign S3[26][2] = S2[26][2];
assign S3[26][3] = S2[26][3];
assign S3[26][4] = S2[26][4];

assign S3[27][0] = S2[27][0];
assign S3[27][1] = S2[27][1];
assign S3[27][2] = S2[27][2];
assign S3[27][3] = S2[27][3];

assign S3[28][0] = S2[28][0];
assign S3[28][1] = S2[28][1];
assign S3[28][2] = S2[28][2];

assign S3[29][0] = S2[29][0];
assign S3[29][1] = S2[29][1];

assign S3[30][0] = S2[30][0];



// S3 - Stage-3 			

assign S4[0][0] = S3[0][0];

assign S4[1][0] = S3[1][0];
assign S4[1][1] = S3[1][1];

assign S4[2][0] = S3[2][0];
assign S4[2][1] = S3[2][1];
assign S4[2][2] = S3[2][2];

assign S4[3][0] = S3[3][0];
assign S4[3][1] = S3[3][1];
assign S4[3][2] = S3[3][2];
assign S4[3][3] = S3[3][3];

assign S4[4][0] = S3[4][0];
assign S4[4][1] = S3[4][1];
assign S4[4][2] = S3[4][2];
assign S4[4][3] = S3[4][3];
assign S4[4][4] = S3[4][4];

assign S4[5][0] = S3[5][0];
assign S4[5][1] = S3[5][1];
assign S4[5][2] = S3[5][2];
assign S4[5][3] = S3[5][3];
assign S4[5][4] = S3[5][4];
assign S4[5][5] = S3[5][5];

HA H301 (S3[6][0], S3[6][1], S4[6][0], S4[7][0]);
assign S4[6][1] = S3[6][2];
assign S4[6][2] = S3[6][3];
assign S4[6][3] = S3[6][4];
assign S4[6][4] = S3[6][5];
assign S4[6][5] = S3[6][6];

FA F301 (S3[7][0], S3[7][1], S3[7][2], S4[7][1], S4[8][0]);
HA H302 (S3[7][3], S3[7][4], S4[7][2], S4[8][1]);
assign S4[7][3] = S3[7][5];
assign S4[7][4] = S3[7][6];
assign S4[7][5] = S3[7][7];

FA F302 (S3[8][0], S3[8][1], S3[8][2], S4[8][2], S4[9][0]);
FA F303 (S3[8][3], S3[8][4], S3[8][5], S4[8][3], S4[9][1]);
HA H303 (S3[8][6], S3[8][7], S4[8][4], S4[9][2]);
assign S4[8][5] = S3[8][8];

genvar k;

generate
	for (k=9; k<=23; k=k+1) begin : block_name_S3
		FA F304 (S3[k][0], S3[k][1], S3[k][2], S4[k][3], S4[k+1][0]);
		FA F305 (S3[k][3], S3[k][4], S3[k][5], S4[k][4], S4[k+1][1]);
		FA F306 (S3[k][6], S3[k][7], S3[k][8], S4[k][5], S4[k+1][2]);
	end

endgenerate


FA F307 (S3[24][0], S3[24][1], S3[24][2], S4[24][3], S4[25][0]);
FA F308 (S3[24][3], S3[24][4], S3[24][5], S4[24][4], S4[25][1]);
assign S4[24][5] = S3[24][6];

FA F309 (S3[25][0], S3[25][1], S3[25][2], S4[25][2], S4[26][0]);
assign S4[25][3] = S3[25][3];
assign S4[25][4] = S3[25][4];
assign S4[25][5] = S3[25][5];

assign S4[26][1] = S3[26][0];
assign S4[26][2] = S3[26][1];
assign S4[26][3] = S3[26][2];
assign S4[26][4] = S3[26][3];
assign S4[26][5] = S3[26][4];

assign S4[27][0] = S3[27][0];
assign S4[27][1] = S3[27][1];
assign S4[27][2] = S3[27][2];
assign S4[27][3] = S3[27][3];

assign S4[28][0] = S3[28][0];
assign S4[28][1] = S3[28][1];
assign S4[28][2] = S3[28][2];

assign S4[29][0] = S3[29][0];
assign S4[29][1] = S3[29][1];

assign S4[30][0] = S3[30][0];




// S4 - Stage-4 			

assign S5[0][0] = S4[0][0];

assign S5[1][0] = S4[1][0];
assign S5[1][1] = S4[1][1];

assign S5[2][0] = S4[2][0];
assign S5[2][1] = S4[2][1];
assign S5[2][2] = S4[2][2];

assign S5[3][0] = S4[3][0];
assign S5[3][1] = S4[3][1];
assign S5[3][2] = S4[3][2];
assign S5[3][3] = S4[3][3];

HA H401 (S4[4][0], S4[4][1], S5[4][0], S5[5][0]);
assign S5[4][1] = S4[4][2];
assign S5[4][2] = S4[4][3];
assign S5[4][3] = S4[4][4];

FA F401 (S4[5][0], S4[5][1], S4[5][2], S5[5][1], S5[6][0]);
HA H402 (S4[5][3], S4[5][4], S5[5][2], S5[6][1]);
assign S5[5][3] = S4[5][5];




genvar k4;

generate

	for(k4=6;k4<=26;k4=k4+1) begin: block_name_S4
		FA F402 (S4[k4][0], S4[k4][1], S4[k4][2], S5[k4][2], S5[k4+1][0]);
		FA F403 (S4[k4][3], S4[k4][4], S4[k4][5], S5[k4][3], S5[k4+1][1]);
	end
	
endgenerate


HA H403 (S4[27][0], S4[27][1], S5[27][2], S5[28][0]);
assign S5[27][3] = S4[27][2];
assign S5[27][4] = S4[27][3];

assign S5[28][1] = S4[28][0];
assign S5[28][2] = S4[28][1];
assign S5[28][3] = S4[28][2];

assign S5[29][0] = S4[29][0];
assign S5[29][1] = S4[29][1];

assign S5[30][0] = S4[30][0];




// S5 - Stage-5 			

assign S6[0][0] = S5[0][0];

assign S6[1][0] = S5[1][0];
assign S6[1][1] = S5[1][1];

assign S6[2][0] = S5[2][0];
assign S6[2][1] = S5[2][1];
assign S6[2][2] = S5[2][2];

HA H501 (S5[3][0], S5[3][1], S6[3][0], S6[4][0]);
assign S6[3][1] = S5[3][2];
assign S6[3][2] = S5[3][3];


genvar k5;

generate

	for(k5=4;k5<=28;k5=k5+1) begin: block_name_S5
		FA F501 (S5[k5][0], S5[k5][1], S5[k5][2], S6[k5][1], S6[k5+1][0]);
		assign S6[k5][2] = S5[k5][3];
	end
	
endgenerate

assign S6[29][1] = S5[29][0];
assign S6[29][2] = S5[29][1];

assign S6[30][0] = S5[30][0];




// S6 - Stage-6 		

assign S7[0][0] = S6[0][0];

assign S7[1][0] = S6[1][0];
assign S7[1][1] = S6[1][1];

HA H601 (S6[2][0], S6[2][1], S7[2][0], S7[3][0]);
assign S7[2][1] = S6[2][2];



genvar k6;

generate

	for(k6=3;k6<=29;k6=k6+1) begin: block_name_S6
		FA F601 (S6[k6][0], S6[k6][1], S6[k6][2], S7[k6][1], S7[k6+1][0]);
	end
	
endgenerate

assign S7[30][1] = S6[30][0];



// RCA

RCA RCA0 ({S7[30][0], S7[29][0], S7[28][0], S7[27][0], S7[26][0], S7[25][0], S7[24][0], S7[23][0], S7[22][0], S7[21][0], S7[20][0], S7[19][0], S7[18][0], S7[17][0], S7[16][0], S7[15][0], S7[14][0], S7[13][0], S7[12][0], S7[11][0], S7[10][0], S7[9][0], S7[8][0], S7[7][0], S7[6][0], S7[5][0], S7[4][0], S7[3][0], S7[2][0], S7[1][0]}, {S7[30][1], S7[29][1], S7[28][1], S7[27][1], S7[26][1], S7[25][1], S7[24][1], S7[23][1], S7[22][1], S7[21][1], S7[20][1], S7[19][1], S7[18][1], S7[17][1], S7[16][1], S7[15][1], S7[14][1], S7[13][1], S7[12][1], S7[11][1], S7[10][1], S7[9][1], S7[8][1], S7[7][1], S7[6][1], S7[5][1], S7[4][1], S7[3][1], S7[2][1], S7[1][1]}, Mul[30:1], Mul[31]);
assign Mul[0] = S7[0][0];

endmodule


module RCA (A, B, Sum, Cout);
input [29:0] A, B;
output Cout;
output [29:0] Sum;

wire C0, C1, C2;

RCA14 R0 (A[13:0], B[13:0], 1'b0, Sum[13:0], C0);
RCA14 R1 (A[27:14], B[27:14], C0, Sum[27:14], C1);
FA F72 (A[28], B[28], C1, Sum[28], C2);
FA F73 (A[29], B[29], C2, Sum[29], Cout);

endmodule


module RCA14 (A, B, Cin, Sum, Cout);
input [13:0] A, B;
input Cin;
output Cout;
output [13:0] Sum;

wire [12:0] C;

FA F59 (A[0], B[0], Cin, Sum[0], C[0]);
FA F60 (A[1], B[1], C[0], Sum[1], C[1]);
FA F61 (A[2], B[2], C[1], Sum[2], C[2]);
FA F62 (A[3], B[3], C[2], Sum[3], C[3]);
FA F63 (A[4], B[4], C[3], Sum[4], C[4]);
FA F64 (A[5], B[5], C[4], Sum[5], C[5]);
FA F65 (A[6], B[6], C[5], Sum[6], C[6]);
FA F66 (A[7], B[7], C[6], Sum[7], C[7]);
FA F67 (A[8], B[8], C[7], Sum[8], C[8]);
FA F68 (A[9], B[9], C[8], Sum[9], C[9]);
FA F69 (A[10], B[10], C[9], Sum[10], C[10]);
FA F70 (A[11], B[11], C[10], Sum[11], C[11]);
FA F71 (A[12], B[12], C[11], Sum[12], C[12]);

FA F72 (A[13], B[13], C[12], Sum[13], Cout);

endmodule




module HA (A, B, Sum, Cout);
input A, B;
output Sum, Cout;

assign Sum = A ^ B;
assign Cout = A & B;

endmodule




module FA(A, B, Cin, Sum, Cout);
input A, B, Cin;
output Sum, Cout;

assign Sum = A ^ B ^ Cin;
assign Cout = ((A ^ B) & Cin) | (A & B);

endmodule
