module Wallace (A, B, Mul);

parameter N = 16;
input [N-1:0] A, B;
output [2*N-1:0] Mul;

reg  S1[31:0][N-1:0];
wire S2[31:0][N-1:0];
wire S3[31:0][N-1:0];
wire S4[31:0][N-1:0];
wire S5[31:0][N-1:0];
wire S6[31:0][N-1:0];
wire S7[31:0][N-1:0];
reg  S8[31:0][N-1:0];

integer i,j,k,m;

always @(*)		// Initialize the partial products (Stage 0)
begin
	for(i=0; i<N; i=i+1)
	begin
		
		for(j=0; j<N; j=j+1)
		begin
			S1[i][j] = A[i] & B[j];
		end
	end
end


// Stage 1				// S stage [weight] [row/# of the element]


assign S2[0][0] = S1[0][0];

HA H1(S1[1][0], S1[0][1], S2[1][0], S2[2][0]);

FA f1 (S1[0][2], S1[1][1], S1[2][0], S2[2][1], S2[3][0]);

FA f2 (S1[0][3], S1[1][2], S1[2][1], S2[3][1], S2[4][0]);
assign S2[3][2] = S1[3][0];

FA f3 (S1[0][4], S1[1][3], S1[2][2], S2[4][1], S2[5][0]);
assign S2[4][2] = S1[3][1];
assign S2[4][3] = S1[4][0];

FA f4 (S1[0][5], S1[1][4], S1[2][3], S2[5][1], S2[6][0]);
FA f5 (S1[3][2], S1[4][1], S1[5][0], S2[5][2], S2[6][1]);

FA f6 (S1[0][6], S1[1][5], S1[2][4], S2[6][2], S2[7][0]);
FA f7 (S1[3][3], S1[4][2], S1[5][1], S2[6][3], S2[7][1]);
assign S2[6][4] = S1[6][0];

FA f8 (S1[0][7], S1[1][6], S1[2][5], S2[7][2], S2[8][0]);
FA f9 (S1[3][4], S1[4][3], S1[5][2], S2[7][3], S2[8][1]);
assign S2[7][4] = S1[6][1];
assign S2[7][5] = S1[7][0];

FA f10 (S1[0][8], S1[1][7], S1[2][6], S2[8][2], S2[9][0]);
FA f11 (S1[3][5], S1[4][4], S1[5][3], S2[8][3], S2[9][1]);
FA f12 (S1[6][2], S1[7][1], S1[8][0], S2[8][4], S2[9][2]);

FA f13 (S1[0][9], S1[1][8], S1[2][7], S2[9][3], S2[10][0]);
FA f14 (S1[3][6], S1[4][5], S1[5][4], S2[9][4], S2[10][1]);
FA f15 (S1[6][3], S1[7][2], S1[8][1], S2[9][5], S2[10][2]);
assign S2[9][6] = S1[9][0];

FA f16 (S1[0][10], S1[1][9], S1[2][8], S2[10][3], S2[11][0]);
FA f17 (S1[3][7] , S1[4][6], S1[5][5], S2[10][4], S2[11][1]);
FA f18 (S1[6][4] , S1[7][3], S1[8][2], S2[10][5], S2[11][2]);
assign S2[10][6] = S1[9][1];
assign S2[10][7] = S1[10][0];

FA f19 (S1[0][11], S1[1][10], S1[2][9] , S2[11][3], S2[12][0]);
FA f20 (S1[3][8] , S1[4][7] , S1[5][6] , S2[11][4], S2[12][1]);
FA f21 (S1[6][5] , S1[7][4] , S1[8][3] , S2[11][5], S2[12][2]);
FA f22 (S1[9][2] , S1[10][1], S1[11][0], S2[11][6], S2[12][3]);

FA f23 (S1[0][12], S1[1][11], S1[2][10], S2[12][4], S2[13][0]);
FA f24 (S1[3][9] , S1[4][8] , S1[5][7] , S2[12][5], S2[13][1]);
FA f25 (S1[6][6] , S1[7][5] , S1[8][4] , S2[12][6], S2[13][2]);
FA f26 (S1[9][3] , S1[10][2], S1[11][1], S2[12][7], S2[13][3]);
assign S2[12][8] = S1[12][0];

FA f27 (S1[0][13], S1[1][12], S1[2][11], S2[13][4], S2[14][0]);
FA f28 (S1[3][10], S1[4][9] , S1[5][8] , S2[13][5], S2[14][1]);
FA f29 (S1[6][7] , S1[7][6] , S1[8][5] , S2[13][6], S2[14][2]);
FA f30 (S1[9][4] , S1[10][3], S1[11][2], S2[13][7], S2[14][3]);
assign S2[13][8] = S1[12][1];
assign S2[13][9] = S1[13][0];

FA f31 (S1[0][14], S1[1][13], S1[2][12], S2[14][4], S2[15][0]);
FA f32 (S1[3][11], S1[4][10], S1[5][9] , S2[14][5], S2[15][1]);
FA f33(S1[6][8] , S1[7][7] , S1[8][6] , S2[14][6], S2[15][2]);
FA f34 (S1[9][5] , S1[10][4], S1[11][3], S2[14][7], S2[15][3]);
FA f35 (S1[12][2], S1[13][1], S1[14][0], S2[14][8], S2[15][4]);

FA f36 (S1[0][15], S1[1][14], S1[2][13], S2[15][5], S2[16][0]);
FA f37 (S1[3][12], S1[4][11], S1[5][10], S2[15][6], S2[16][1]);
FA f38 (S1[6][9] , S1[7][8] , S1[8][7] , S2[15][7], S2[16][2]);
FA f39 (S1[9][6] , S1[10][5], S1[11][4], S2[15][8], S2[16][3]);
FA f40 (S1[12][3], S1[13][2], S1[14][1], S2[15][9], S2[16][4]);
assign S2[15][10] = S1[15][0];

FA f41 (S1[15][1], S1[14][2], S1[13][3], S2[16][5], S2[17][0]);
FA f42 (S1[12][4], S1[11][5], S1[10][6], S2[16][6], S2[17][1]);
FA f43 (S1[9][7] , S1[8][8] , S1[7][9] , S2[16][7], S2[17][2]);
FA f44 (S1[6][10], S1[5][11], S1[4][12], S2[16][8], S2[17][3]);
FA f45 (S1[3][13], S1[2][14], S1[1][15], S2[16][9], S2[17][4]);

FA f46 (S1[15][2], S1[14][3], S1[13][4], S2[17][5], S2[18][0]);
FA f47 (S1[12][5], S1[11][6], S1[10][7], S2[17][6], S2[18][1]);
FA f48 (S1[9][8] , S1[8][9] , S1[7][10], S2[17][7], S2[18][2]);
FA f49 (S1[6][11], S1[5][12], S1[4][13], S2[17][8], S2[18][3]);
assign S2[17][9]  = S1[3][14];
assign S2[17][10] = S1[2][15];

FA f50 (S1[15][3], S1[14][4], S1[13][5], S2[18][4], S2[19][0]);
FA f51 (S1[12][6], S1[11][7], S1[10][8], S2[18][5], S2[19][1]);
FA f52 (S1[9][9] , S1[8][10], S1[7][11], S2[18][6], S2[19][2]);
FA f53 (S1[6][12], S1[5][13], S1[4][14], S2[18][7], S2[19][3]);
assign S2[18][8] = S1[3][15];

FA f54 (S1[15][4], S1[14][5], S1[13][6], S2[19][4], S2[20][0]);
FA f55(S1[12][7], S1[11][8], S1[10][9], S2[19][5], S2[20][1]);
FA f56 (S1[9][10], S1[8][11], S1[7][12], S2[19][6], S2[20][2]);
FA f57 (S1[6][13], S1[5][14], S1[4][15], S2[19][7], S2[20][3]);

FA f58 (S1[15][5], S1[14][6], S1[13][7] , S2[20][4], S2[21][0]);
FA f59 (S1[12][8], S1[11][9], S1[10][10], S2[20][5], S2[21][1]);
FA f60 (S1[9][11], S1[8][12], S1[7][13] , S2[20][6], S2[21][2]);
assign S2[20][7] = S1[6][14];
assign S2[20][8] = S1[5][15];

FA f61 (S1[15][6], S1[14][7] , S1[13][8] , S2[21][3], S2[22][0]);
FA f62 (S1[12][9], S1[11][10], S1[10][11], S2[21][4], S2[22][1]);
FA f63 (S1[9][12], S1[8][13] , S1[7][14] , S2[21][5], S2[22][2]);
assign S2[21][6] = S1[6][15];

FA f64 (S1[15][7] , S1[14][8] , S1[13][9] , S2[22][3], S2[23][0]);
FA f65 (S1[12][10], S1[11][11], S1[10][12], S2[22][4], S2[23][1]);
FA f66 (S1[9][13] , S1[8][14] , S1[7][15] , S2[22][5], S2[23][2]);

FA f67 (S1[15][8] , S1[14][9] , S1[13][10], S2[23][3], S2[24][0]);
FA f68 (S1[12][11], S1[11][12], S1[10][13], S2[23][4], S2[24][1]);
assign S2[23][5] = S1[9][14];
assign S2[23][6] = S1[8][15];

FA f69 (S1[15][9] , S1[14][10], S1[13][11], S2[24][2], S2[25][0]);
FA f70 (S1[12][12], S1[11][13], S1[10][14], S2[24][3], S2[25][1]);
assign S2[24][4] = S1[9][15];

FA f71 (S1[15][10], S1[14][11], S1[13][12], S2[25][2], S2[26][0]);
FA f72 (S1[12][13], S1[11][14], S1[10][15], S2[25][3], S2[26][1]);

FA f73 (S1[15][11], S1[14][12], S1[13][13], S2[26][2], S2[27][0]);
assign S2[26][3] = S1[12][14];
assign S2[26][4] = S1[11][15];

FA f74 (S1[15][12], S1[14][13], S1[13][14], S2[27][1], S2[28][0]);
assign S2[27][2] = S1[12][15];

FA f75 (S1[15][13], S1[14][14], S1[13][15], S2[28][1], S2[29][0]);

assign S2[29][1] = S1[15][14];
assign S2[29][2] = S1[14][15];

assign S2[30][0] = S1[15][15];




// Stage 2				// S stage [weight] [row/# of the element]

assign S3[0][0] = S2[0][0];

assign S3[1][0] = S2[1][0];

HA H2 (S2[2][0], S2[2][1], S3[2][0], S3[3][0]);

FA f101 (S2[3][0], S2[3][1], S2[3][2], S3[3][1], S3[4][0]);

FA f102 (S2[4][0], S2[4][1], S2[4][2], S3[4][1], S3[5][0]);
assign S3[4][2] = S2[4][3];

FA f103(S2[5][0], S2[5][1], S2[5][2], S3[5][1], S3[6][0]);

FA f104 (S2[6][0], S2[6][1], S2[6][2], S3[6][1], S3[7][0]);
assign S3[6][2] = S2[6][3];
assign S3[6][3] = S2[6][4];

FA f105 (S2[7][0], S2[7][1], S2[7][2], S3[7][1], S3[8][0]);
FA f106 (S2[7][3], S2[7][4], S2[7][5], S3[7][2], S3[8][1]);

FA f107 (S2[8][0], S2[8][1], S2[8][2], S3[8][2], S3[9][0]);
assign S3[8][3] = S2[8][3];
assign S3[8][4] = S2[8][4];

FA f108 (S2[9][0], S2[9][1], S2[9][2], S3[9][1], S3[10][0]);
FA f109 (S2[9][3], S2[9][4], S2[9][5], S3[9][2], S3[10][1]);
assign S3[9][3] = S2[9][6]; 

FA f110 (S2[10][0], S2[10][1], S2[10][2], S3[10][2], S3[11][0]);
FA f111 (S2[10][3], S2[10][4], S2[10][5], S3[10][3], S3[11][1]);
assign S3[10][4] = S2[10][6];
assign S3[10][5] = S2[10][7];

FA f112 (S2[11][0], S2[11][1], S2[11][2], S3[11][2], S3[12][0]);
FA f113(S2[11][3], S2[11][4], S2[11][5], S3[11][3], S3[12][1]);
assign S3[11][4] = S2[11][6];

FA f114 (S2[12][0], S2[12][1], S2[12][2], S3[12][2], S3[13][0]);
FA f115 (S2[12][3], S2[12][4], S2[12][5], S3[12][3], S3[13][1]);
FA f116 (S2[12][6], S2[12][7], S2[12][8], S3[12][4], S3[13][2]);

FA f117 (S2[13][0], S2[13][1], S2[13][2], S3[13][3], S3[14][0]);
FA f118 (S2[13][3], S2[13][4], S2[13][5], S3[13][4], S3[14][1]);
FA f119 (S2[13][6], S2[13][7], S2[13][8], S3[13][5], S3[14][2]);
assign S3[13][6] = S2[13][9];

FA f120 (S2[14][0], S2[14][1], S2[14][2], S3[14][3], S3[15][0]);
FA f121 (S2[14][3], S2[14][4], S2[14][5], S3[14][4], S3[15][1]);
FA f122 (S2[14][6], S2[14][7], S2[14][8], S3[14][5], S3[15][2]);

FA f123 (S2[15][0], S2[15][1], S2[15][2], S3[15][3], S3[16][0]);
FA f124 (S2[15][3], S2[15][4], S2[15][5], S3[15][4], S3[16][1]);
FA f125 (S2[15][6], S2[15][7], S2[15][8], S3[15][5], S3[16][2]);
assign S3[15][6] = S2[15][9] ;
assign S3[15][7] = S2[15][10];

FA f126 (S2[16][0], S2[16][1], S2[16][2], S3[16][3], S3[17][0]);
FA f127 (S2[16][3], S2[16][4], S2[16][5], S3[16][4], S3[17][1]);
FA f128 (S2[16][6], S2[16][7], S2[16][8], S3[16][5], S3[17][2]);
assign S3[16][6] = S2[16][9] ;

FA f129 (S2[17][0], S2[17][1], S2[17][2], S3[17][3], S3[18][0]);
FA f130 (S2[17][3], S2[17][4], S2[17][5], S3[17][4], S3[18][1]);
FA f131 (S2[17][6], S2[17][7], S2[17][8], S3[17][5], S3[18][2]);
assign S3[17][6] = S2[17][9] ;
assign S3[17][7] = S2[17][10];

FA f132 (S2[18][0], S2[18][1], S2[18][2], S3[18][3], S3[19][0]);
FA f133 (S2[18][3], S2[18][4], S2[18][5], S3[18][4], S3[19][1]);
FA f134 (S2[18][6], S2[18][7], S2[18][8], S3[18][5], S3[19][2]);

FA f135 (S2[19][0], S2[19][1], S2[19][2], S3[19][3], S3[20][0]);
FA f136 (S2[19][3], S2[19][4], S2[19][5], S3[19][4], S3[20][1]);
assign S3[19][5] = S2[19][6];
assign S3[19][6] = S2[19][7];

FA f137 (S2[20][0], S2[20][1], S2[20][2], S3[20][2], S3[21][0]);
FA f138 (S2[20][3], S2[20][4], S2[20][5], S3[20][3], S3[21][1]);
FA f139 (S2[20][6], S2[20][7], S2[20][8], S3[20][4], S3[21][2]);

FA f140 (S2[21][0], S2[21][1], S2[21][2], S3[21][3], S3[22][0]);
FA f141 (S2[21][3], S2[21][4], S2[21][5], S3[21][4], S3[22][1]);
assign S3[21][5] = S2[21][6];

FA f142 (S2[22][0], S2[22][1], S2[22][2], S3[22][2], S3[23][0]);
FA f143 (S2[22][3], S2[22][4], S2[22][5], S3[22][3], S3[23][1]);

FA f144 (S2[23][0], S2[23][1], S2[23][2], S3[23][2], S3[24][0]);
FA f145 (S2[23][3], S2[23][4], S2[23][5], S3[23][3], S3[24][1]);
assign S3[23][4] = S2[23][6];

FA f146 (S2[24][0], S2[24][1], S2[24][2], S3[24][2], S3[25][0]);
assign S3[24][3] = S2[24][3];
assign S3[24][4] = S2[24][4];

FA f147 (S2[25][0], S2[25][1], S2[25][2], S3[25][1], S3[26][0]);
assign S3[25][2] = S2[25][3];

FA f148 (S2[26][0], S2[26][1], S2[26][2], S3[26][1], S3[27][0]);
assign S3[26][2] = S2[26][3];
assign S3[26][3] = S2[26][4];

FA f149 (S2[27][0], S2[27][1], S2[27][2], S3[27][1], S3[28][0]);

assign S3[28][1] = S2[28][0];
assign S3[28][2] = S2[28][1];

FA f150 (S2[29][0], S2[29][1], S2[29][2], S3[29][0], S3[30][0]);

assign S3[30][1] = S2[30][0];




// Stage 3				// S stage [weight] [row/# of the element]

assign S4[0][0] = S3[0][0];

assign S4[1][0] = S3[1][0];

assign S4[2][0] = S3[2][0];

HA H3 (S3[3][0], S3[3][1], S4[3][0], S4[4][0]);

FA f201 (S3[4][0], S3[4][1], S3[4][2], S4[4][1], S4[5][0]);

assign S4[5][1] = S3[5][0];
assign S4[5][2] = S3[5][1];

FA f202 (S3[6][0], S3[6][1], S3[6][2], S4[6][0], S4[7][0]);
assign S4[6][1] = S3[6][3];

FA f203 (S3[7][0], S3[7][1], S3[7][2], S4[7][1], S4[8][0]);

FA f204 (S3[8][0], S3[8][1], S3[8][2], S4[8][1], S4[9][0]);
assign S4[8][2] = S3[8][3];
assign S4[8][3] = S3[8][4];

FA f205 (S3[9][0], S3[9][1], S3[9][2], S4[9][1], S4[10][0]);
assign S4[9][2] = S3[9][3];

FA f206 (S3[10][0], S3[10][1], S3[10][2], S4[10][1], S4[11][0]);
FA f207 (S3[10][3], S3[10][4], S3[10][5], S4[10][2], S4[11][1]);

FA f208 (S3[11][0], S3[11][1], S3[11][2], S4[11][2], S4[12][0]);
assign S4[11][3] = S3[11][3];
assign S4[11][4] = S3[11][4];

FA f209 (S3[12][0], S3[12][1], S3[12][2], S4[12][1], S4[13][0]);
assign S4[12][2] = S3[12][3];
assign S4[12][3] = S3[12][4];

FA f210 (S3[13][0], S3[13][1], S3[13][2], S4[13][1], S4[14][0]);
FA f211 (S3[13][3], S3[13][4], S3[13][5], S4[13][2], S4[14][1]);
assign S4[13][3] = S3[13][6];

FA f212 (S3[14][0], S3[14][1], S3[14][2], S4[14][2], S4[15][0]);
FA f213 (S3[14][3], S3[14][4], S3[14][5], S4[14][3], S4[15][1]);

FA f214 (S3[15][0], S3[15][1], S3[15][2], S4[15][2], S4[16][0]);
FA f215 (S3[15][3], S3[15][4], S3[15][5], S4[15][3], S4[16][1]);
assign S4[15][4] = S3[15][6];
assign S4[15][5] = S3[15][7];

FA f216 (S3[16][0], S3[16][1], S3[16][2], S4[16][2], S4[17][0]);
FA f217 (S3[16][3], S3[16][4], S3[16][5], S4[16][3], S4[17][1]);
assign S4[16][4] = S3[16][6];

FA f218 (S3[17][0], S3[17][1], S3[17][2], S4[17][2], S4[18][0]);
FA f219 (S3[17][3], S3[17][4], S3[17][5], S4[17][3], S4[18][1]);
assign S4[17][4] = S3[17][6];
assign S4[17][5] = S3[17][7];

FA f220 (S3[18][0], S3[18][1], S3[18][2], S4[18][2], S4[19][0]);
FA f221 (S3[18][3], S3[18][4], S3[18][5], S4[18][3], S4[19][1]);

FA f222 (S3[19][0], S3[19][1], S3[19][2], S4[19][2], S4[20][0]);
FA f223 (S3[19][3], S3[19][4], S3[19][5], S4[19][3], S4[20][1]);
assign S4[19][4] = S3[19][6];

FA f224 (S3[20][0], S3[20][1], S3[20][2], S4[20][2], S4[21][0]);
assign S4[20][3] = S3[20][3];
assign S4[20][4] = S3[20][4];

FA f225 (S3[21][0], S3[21][1], S3[21][2], S4[21][1], S4[22][0]);
FA f226 (S3[21][3], S3[21][4], S3[21][5], S4[21][2], S4[22][1]);

FA f227 (S3[22][0], S3[22][1], S3[22][2], S4[22][2], S4[23][0]);
assign S4[22][3] = S3[22][3];

FA f228 (S3[23][0], S3[23][1], S3[23][2], S4[23][1], S4[24][0]);
assign S4[23][2] = S3[23][3];
assign S4[23][3] = S3[23][4];

FA f229 (S3[24][0], S3[24][1], S3[24][2], S4[24][1], S4[25][0]);
assign S4[24][2] = S3[24][3];
assign S4[24][3] = S3[24][4];

FA f230 (S3[25][0], S3[25][1], S3[25][2], S4[25][1], S4[26][0]);

FA f231 (S3[26][0], S3[26][1], S3[26][2], S4[26][1], S4[27][0]);
assign S4[26][2] = S3[26][3];

assign S4[27][1] = S3[27][0];
assign S4[27][2] = S3[27][1];

FA f232 (S3[28][0], S3[28][1], S3[28][2], S4[28][0], S4[29][0]);

assign S4[29][1] = S3[29][0];

assign S4[30][0] = S3[30][0];
assign S4[30][1] = S3[30][1];



// Stage 4				// S stage [weight] [row/# of the element]

assign S5[0][0] = S4[0][0];

assign S5[1][0] = S4[1][0];

assign S5[2][0] = S4[2][0];

assign S5[3][0] = S4[3][0];

HA H4 (S4[4][0], S4[4][1], S5[4][0], S5[5][0]);

FA f301 (S4[5][0], S4[5][1], S4[5][2], S5[5][1], S5[6][0]);

assign S5[6][1] = S4[6][0];
assign S5[6][2] = S4[6][1];

assign S5[7][0] = S4[7][0];
assign S5[7][1] = S4[7][1];

FA f302 (S4[8][0], S4[8][1], S4[8][2], S5[8][0], S5[9][0]);
assign S5[8][1] = S4[8][3];

FA f303 (S4[9][0], S4[9][1], S4[9][2], S5[9][1], S5[10][0]);

FA f304 (S4[10][0], S4[10][1], S4[10][2], S5[10][1], S5[11][0]);

FA f305 (S4[11][0], S4[11][1], S4[11][2], S5[11][1], S5[12][0]);
assign S5[11][2] = S4[11][3];
assign S5[11][3] = S4[11][4];

FA f306 (S4[12][0], S4[12][1], S4[12][2], S5[12][1], S5[13][0]);
assign S5[12][2] = S4[12][3];

FA f307 (S4[13][0], S4[13][1], S4[13][2], S5[13][1], S5[14][0]);
assign S5[13][2] = S4[13][3];

FA f308 (S4[14][0], S4[14][1], S4[14][2], S5[14][1], S5[15][0]);
assign S5[14][2] = S4[14][3];

FA f309 (S4[15][0], S4[15][1], S4[15][2], S5[15][1], S5[16][0]);
FA f310 (S4[15][3], S4[15][4], S4[15][5], S5[15][2], S5[16][1]);

FA f311 (S4[16][0], S4[16][1], S4[16][2], S5[16][2], S5[17][0]);
HA H5 (S4[16][3], S4[16][4], S5[16][3], S5[17][1]);

FA f312 (S4[17][0], S4[17][1], S4[17][2], S5[17][2], S5[18][0]);
FA f313 (S4[17][3], S4[17][4], S4[17][5], S5[17][3], S5[18][1]);

FA f314 (S4[18][0], S4[18][1], S4[18][2], S5[18][2], S5[19][0]);
assign S5[18][3] = S4[18][3];

FA f315 (S4[19][0], S4[19][1], S4[19][2], S5[19][1], S5[20][0]);
assign S5[19][2] = S4[19][3];
assign S5[19][3] = S4[19][4];

FA f316 (S4[20][0], S4[20][1], S4[20][2], S5[20][1], S5[21][0]);
assign S5[20][2] = S4[20][3];
assign S5[20][3] = S4[20][4];

FA f317 (S4[21][0], S4[21][1], S4[21][2], S5[21][1], S5[22][0]);

FA f318 (S4[22][0], S4[22][1], S4[22][2], S5[22][1], S5[23][0]);
assign S5[22][2] = S4[22][3];

FA f319 (S4[23][0], S4[23][1], S4[23][2], S5[23][1], S5[24][0]);
assign S5[23][2] = S4[23][3];

FA f320 (S4[24][0], S4[24][1], S4[24][2], S5[24][1], S5[25][0]);
assign S5[24][2] = S4[24][3];

assign S5[25][1] = S4[25][0];
assign S5[25][2] = S4[25][1];

FA f321 (S4[26][0], S4[26][1], S4[26][2], S5[26][0], S5[27][0]);

FA f322 (S4[27][0], S4[27][1], S4[27][2], S5[27][1], S5[28][0]);

assign S5[28][1] = S4[28][0];

assign S5[29][0] = S4[29][0];
assign S5[29][1] = S4[29][1];

assign S5[30][0] = S4[30][0];
assign S5[30][1] = S4[30][1];



// Stage 5				// S stage [weight] [row/# of the element]

assign S6[0][0] = S5[0][0];

assign S6[1][0] = S5[1][0];

assign S6[2][0] = S5[2][0];

assign S6[3][0] = S5[3][0];

assign S6[4][0] = S5[4][0];

HA H15 (S5[5][0], S5[5][1], S6[5][0], S6[6][0]);

FA f401 (S5[6][0], S5[6][1], S5[6][2], S6[6][1], S6[7][0]);

assign S6[7][1] = S5[7][0];
assign S6[7][2] = S5[7][1];

assign S6[8][0] = S5[8][0];
assign S6[8][1] = S5[8][1];

assign S6[9][0] = S5[9][0];
assign S6[9][1] = S5[9][1];

assign S6[10][0] = S5[10][0];
assign S6[10][1] = S5[10][1];

FA f402 (S5[11][0], S5[11][1], S5[11][2], S6[11][0], S6[12][0]);
assign S6[11][1] = S5[11][3];

FA f403 (S5[12][0], S5[12][1], S5[12][2], S6[12][1], S6[13][0]);

FA f404 (S5[13][0], S5[13][1], S5[13][2], S6[13][1], S6[14][0]);

FA f405 (S5[14][0], S5[14][1], S5[14][2], S6[14][1], S6[15][0]);

FA f406 (S5[15][0], S5[15][1], S5[15][2], S6[15][1], S6[16][0]);

FA f407 (S5[16][0], S5[16][1], S5[16][2], S6[16][1], S6[17][0]);
assign S6[16][2] = S5[16][3];

FA f408 (S5[17][0], S5[17][1], S5[17][2], S6[17][1], S6[18][0]);
assign S6[17][2] = S5[17][3];

FA f409 (S5[18][0], S5[18][1], S5[18][2], S6[18][1], S6[19][0]);
assign S6[18][2] = S5[18][3];

FA f410 (S5[19][0], S5[19][1], S5[19][2], S6[19][1], S6[20][0]);
assign S6[19][2] = S5[19][3];

FA f411 (S5[20][0], S5[20][1], S5[20][2], S6[20][1], S6[21][0]);
assign S6[20][2] = S5[20][3];

assign S6[21][1] = S5[21][0];
assign S6[21][2] = S5[21][1];

FA f412 (S5[22][0], S5[22][1], S5[22][2], S6[22][0], S6[23][0]);

FA f413 (S5[23][0], S5[23][1], S5[23][2], S6[23][1], S6[24][0]);

FA f414 (S5[24][0], S5[24][1], S5[24][2], S6[24][1], S6[25][0]);

FA f415 (S5[25][0], S5[25][1], S5[25][2], S6[25][1], S6[26][0]);

assign S6[26][1] = S5[26][0];

assign S6[27][0] = S5[27][0];
assign S6[27][1] = S5[27][1];

assign S6[28][0] = S5[28][0];
assign S6[28][1] = S5[28][1];

assign S6[29][0] = S5[29][0];
assign S6[29][1] = S5[29][1];

assign S6[30][0] = S5[30][0];
assign S6[30][1] = S5[30][1];



// Stage 5				// S stage [weight] [row/# of the element]

assign S7[0][0] = S6[0][0];

assign S7[1][0] = S6[1][0];

assign S7[2][0] = S6[2][0];

assign S7[3][0] = S6[3][0];

assign S7[4][0] = S6[4][0];

assign S7[5][0] = S6[5][0];

HA H6 (S6[6][0], S6[6][1], S7[6][0], S7[7][0]);

FA f501 (S6[7][0], S6[7][1], S6[7][2], S7[7][1], S7[8][0]);

HA H7 (S6[8][0], S6[8][1], S7[8][1], S7[9][0]);

HA H8 (S6[9][0], S6[9][1], S7[9][1], S7[10][0]);

HA H9 (S6[10][0], S6[10][1], S7[10][1], S7[11][0]);

HA H10 (S6[11][0], S6[11][1], S7[11][1], S7[12][0]);

HA H11 (S6[12][0], S6[12][1], S7[12][1], S7[13][0]);

HA H12 (S6[13][0], S6[13][1], S7[13][1], S7[14][0]);

HA H13 (S6[14][0], S6[14][1], S7[14][1], S7[15][0]);

HA H14 (S6[15][0], S6[15][1], S7[15][1], S7[16][0]);

FA f502 (S6[16][0], S6[16][1], S6[16][2], S7[16][1], S7[17][0]);

FA f503 (S6[17][0], S6[17][1], S6[17][2], S7[17][1], S7[18][0]);

FA f504 (S6[18][0], S6[18][1], S6[18][2], S7[18][1], S7[19][0]);

FA f505 (S6[19][0], S6[19][1], S6[19][2], S7[19][1], S7[20][0]);

FA f506 (S6[20][0], S6[20][1], S6[20][2], S7[20][1], S7[21][0]);

FA f507 (S6[21][0], S6[21][1], S6[21][2], S7[21][1], S7[22][0]);

assign S7[22][1] = S6[22][0];

assign S7[23][0] = S6[23][0];
assign S7[23][1] = S6[23][1];

assign S7[24][0] = S6[24][0];
assign S7[24][1] = S6[24][1];

assign S7[25][0] = S6[25][0];
assign S7[25][1] = S6[25][1];

assign S7[26][0] = S6[26][0];
assign S7[26][1] = S6[26][1];

assign S7[27][0] = S6[27][0];
assign S7[27][1] = S6[27][1];

assign S7[28][0] = S6[28][0];
assign S7[28][1] = S6[28][1];

assign S7[29][0] = S6[29][0];
assign S7[29][1] = S6[29][1];

assign S7[30][0] = S6[30][0];
assign S7[30][1] = S6[30][1];



// Stage 6				// S stage [weight] [row/# of the element]


// assign S8[0][0] = S7[0][0];

// assign S8[1][0] = S7[1][0];

// assign S8[2][0] = S7[2][0];

// assign S8[3][0] = S7[3][0];

// assign S8[4][0] = S7[4][0];

// assign S8[5][0] = S7[5][0];

// assign S8[6][0] = S7[6][0];


always @(*)
begin
	for (k=0;k<7;k=k+1)
		S8[k][0] = S7[k][0];
end



// assign S8[7][0] = S7[7][0];
// assign S8[7][1] = S7[7][1];

always @(*) begin
	for (m=7;m<31;m=m+1)
	begin
		S8[m][0] = S7[m][0];
		S8[m][1] = S7[m][1];
	end
end


assign Mul[6:0] = {S8[6][0], S8[5][0], S8[4][0], S8[3][0], S8[2][0], S8[1][0], S8[0][0]};
// 24-bit Ripple Carry Adder

RCA24 RC0 ({S8[30][0], S8[29][0], S8[28][0], S8[27][0], S8[26][0], S8[25][0], S8[24][0], S8[23][0], S8[22][0], S8[21][0], S8[20][0], S8[19][0], S8[18][0], S8[17][0], S8[16][0], S8[15][0], S8[14][0], S8[13][0], S8[12][0], S8[11][0], S8[10][0], S8[9][0], S8[8][0], S8[7][0]}, {S8[30][1], S8[29][1], S8[28][1], S8[27][1], S8[26][1], S8[25][1], S8[24][1], S8[23][1], S8[22][1], S8[21][1], S8[20][1], S8[19][1], S8[18][1], S8[17][1], S8[16][1], S8[15][1], S8[14][1], S8[13][1], S8[12][1], S8[11][1], S8[10][1], S8[9][1], S8[8][1], S8[7][1]}, Mul[30:7], Mul[31]);


endmodule


// 24-bit RCA

module RCA24 (A, B, Sum, Cout);
input [23:0] A, B;
output [23:0] Sum;
output Cout;
wire C;

RCA12 R1 (A[11:0] , B[11:0] , 1'b0, Sum[11:0] , C);
RCA12 R2 (A[23:12], B[23:12], C,    Sum[23:12], Cout);

endmodule

module RCA12 (A, B, Cin, Sum, Cout);
input [11:0] A, B;
input Cin;
output Cout;
output [11:0] Sum;

wire [10:0] C;

FA H959 (A[0], B[0], Cin , Sum[0], C[0]);
FA F960 (A[1], B[1], C[0], Sum[1], C[1]);
FA F961 (A[2], B[2], C[1], Sum[2], C[2]);
FA F962 (A[3], B[3], C[2], Sum[3], C[3]);
FA F963 (A[4], B[4], C[3], Sum[4], C[4]);
FA F964 (A[5], B[5], C[4], Sum[5], C[5]);
FA F965 (A[6], B[6], C[5], Sum[6], C[6]);
FA F966 (A[7], B[7], C[6], Sum[7], C[7]);
FA F967 (A[8], B[8], C[7], Sum[8], C[8]);
FA F968 (A[9], B[9], C[8], Sum[9], C[9]);

FA F969 (A[10], B[10], C[9] , Sum[10], C[10]);
FA F970 (A[11], B[11], C[10], Sum[11], Cout );
endmodule



// Half_Adder

module HA (A, B, Sum, Cout);
input A, B;
output Sum, Cout;

assign Sum = A ^ B;
assign Cout = A & B;

endmodule


// Full_Adder

module FA(A, B, Cin, Sum, Cout);
input A, B, Cin;
output Sum, Cout;

assign Sum = A ^ B ^ Cin;
assign Cout = ((A ^ B) & Cin) | (A & B);

endmodule